`timescale 1 ps / 1 ps

/***
*
*	task2RAM module
* 	builds a 32x3 memory file using a memory array
* 	takes in 5bit address, to be read and written to
*	takes in 3 bit data in, for data to be written
* 	takes in 1 bit CLOCK_50 and wren, for clock and write enable
* 	outputs 3 bit q, for data out
*
*
***/
module task2RAM (	address, CLOCK_50, data, wren, q);
	input	logic [4:0]  address;
	input	logic 		 CLOCK_50;
	input	logic [2:0]  data;
	input	logic 		 wren;
	output logic [2:0]  q;
	
	assign clock = CLOCK_50;
	
	logic [2:0] memory_array [31:0];
	
	always_ff @(posedge clock) begin
		if(wren) begin
			memory_array[address] <= data;
			q <= data;
		
		end else begin
			q <= memory_array[address];
		end	
	
	end
	
endmodule

module task2RAM_testbench ();
	logic	[4:0]  address;
	logic	  		 clock;
	logic	[2:0]  data;
	logic	  		 wren;
	logic [2:0]  q;
	
	task2RAM dut (.address(address), .CLOCK_50(clock), .data(data), .wren(wren), .q(q));

	 // Set up a simulated clock.   
	parameter CLOCK_PERIOD=100; 

	initial begin   
		clock <= 0;  
		forever #(CLOCK_PERIOD/2) clock <= ~clock; // Forever toggle the clock 
	end  
		
	// Test the design. 
	initial begin  
																	   @(posedge clock);
	wren <= 0;  address [4:0] <= 0;  data [2:0] <= 0;  @(posedge clock); // set all values to 0
												data [0] <= 1;		@(posedge clock); // cycling through all 8 variations of bit representation
						   data [1] <= 1; data [0] <= 0;		@(posedge clock);
												data [0] <= 1;		@(posedge clock);
							data [2] <= 1;	data [1:0] <= 0;  @(posedge clock);
												data [0] <= 1;		@(posedge clock);
						   data [1] <= 1; data [0] <= 0;		@(posedge clock);
												data [0] <= 1;		@(posedge clock);
							data [3] <= 1; data [2:0] <= 0;  @(posedge clock);
												data [0] <= 1;		@(posedge clock);
						   data [1] <= 1; data [0] <= 0;		@(posedge clock);
												data [0] <= 1;		@(posedge clock);
							data [2] <= 1;	data [1:0] <= 0;  @(posedge clock);
												data [0] <= 1;		@(posedge clock);
						   data [1] <= 1; data [0] <= 0;		@(posedge clock);
												data [0] <= 1;		@(posedge clock);
					address [0] <= 1;								@(posedge clock); // through 32 variations of bit representation
							data [0] <= 1;							@(posedge clock); // each address bit representation cycles through
						   data [1] <= 1; data [0] <= 0;		@(posedge clock); // all 8 variations of data representation
												data [0] <= 1;		@(posedge clock);
							data [2] <= 1;	data [1:0] <= 0;  @(posedge clock);
												data [0] <= 1;		@(posedge clock);
						   data [1] <= 1; data [0] <= 0;		@(posedge clock);
												data [0] <= 1;		@(posedge clock);
							data [3] <= 1; data [2:0] <= 0;  @(posedge clock);
												data [0] <= 1;		@(posedge clock);
						   data [1] <= 1; data [0] <= 0;		@(posedge clock);
												data [0] <= 1;		@(posedge clock);
							data [2] <= 1;	data [1:0] <= 0;  @(posedge clock);
												data [0] <= 1;		@(posedge clock);
						   data [1] <= 1; data [0] <= 0;		@(posedge clock);
												data [0] <= 1;		@(posedge clock);
					address [1] <= 1; address [0] <= 0;		@(posedge clock);
							data [0] <= 1;							@(posedge clock);
						   data [1] <= 1; data [0] <= 0;		@(posedge clock);
												data [0] <= 1;		@(posedge clock);
							data [2] <= 1;	data [1:0] <= 0;  @(posedge clock);
												data [0] <= 1;		@(posedge clock);
						   data [1] <= 1; data [0] <= 0;		@(posedge clock);
												data [0] <= 1;		@(posedge clock);
							data [3] <= 1; data [2:0] <= 0;  @(posedge clock);
												data [0] <= 1;		@(posedge clock);
						   data [1] <= 1; data [0] <= 0;		@(posedge clock);
												data [0] <= 1;		@(posedge clock);
							data [2] <= 1;	data [1:0] <= 0;  @(posedge clock);
												data [0] <= 1;		@(posedge clock);
						   data [1] <= 1; data [0] <= 0;		@(posedge clock);
												data [0] <= 1;		@(posedge clock);					
					address [0] <= 1;								@(posedge clock);
							data [0] <= 1;							@(posedge clock);
						   data [1] <= 1; data [0] <= 0;		@(posedge clock);
												data [0] <= 1;		@(posedge clock);
							data [2] <= 1;	data [1:0] <= 0;  @(posedge clock);
												data [0] <= 1;		@(posedge clock);
						   data [1] <= 1; data [0] <= 0;		@(posedge clock);
												data [0] <= 1;		@(posedge clock);
							data [3] <= 1; data [2:0] <= 0;  @(posedge clock);
												data [0] <= 1;		@(posedge clock);
						   data [1] <= 1; data [0] <= 0;		@(posedge clock);
												data [0] <= 1;		@(posedge clock);
							data [2] <= 1;	data [1:0] <= 0;  @(posedge clock);
												data [0] <= 1;		@(posedge clock);
						   data [1] <= 1; data [0] <= 0;		@(posedge clock);
												data [0] <= 1;		@(posedge clock);					
					address [2] <= 1; address [1:0] <= 0;  @(posedge clock);
							data [0] <= 1;							@(posedge clock);
						   data [1] <= 1; data [0] <= 0;		@(posedge clock);
												data [0] <= 1;		@(posedge clock);
							data [2] <= 1;	data [1:0] <= 0;  @(posedge clock);
												data [0] <= 1;		@(posedge clock);
						   data [1] <= 1; data [0] <= 0;		@(posedge clock);
												data [0] <= 1;		@(posedge clock);
							data [3] <= 1; data [2:0] <= 0;  @(posedge clock);
												data [0] <= 1;		@(posedge clock);
						   data [1] <= 1; data [0] <= 0;		@(posedge clock);
												data [0] <= 1;		@(posedge clock);
							data [2] <= 1;	data [1:0] <= 0;  @(posedge clock);
												data [0] <= 1;		@(posedge clock);
						   data [1] <= 1; data [0] <= 0;		@(posedge clock);
												data [0] <= 1;		@(posedge clock);					
					address [0] <= 1; 							@(posedge clock);
							data [0] <= 1;							@(posedge clock);
						   data [1] <= 1; data [0] <= 0;		@(posedge clock);
												data [0] <= 1;		@(posedge clock);
							data [2] <= 1;	data [1:0] <= 0;  @(posedge clock);
												data [0] <= 1;		@(posedge clock);
						   data [1] <= 1; data [0] <= 0;		@(posedge clock);
												data [0] <= 1;		@(posedge clock);
							data [3] <= 1; data [2:0] <= 0;  @(posedge clock);
												data [0] <= 1;		@(posedge clock);
						   data [1] <= 1; data [0] <= 0;		@(posedge clock);
												data [0] <= 1;		@(posedge clock);
							data [2] <= 1;	data [1:0] <= 0;  @(posedge clock);
												data [0] <= 1;		@(posedge clock);
						   data [1] <= 1; data [0] <= 0;		@(posedge clock);
												data [0] <= 1;		@(posedge clock);					
					address [1] <= 1; address [0] <= 0;    @(posedge clock);
							data [0] <= 1;							@(posedge clock);
						   data [1] <= 1; data [0] <= 0;		@(posedge clock);
												data [0] <= 1;		@(posedge clock);
							data [2] <= 1;	data [1:0] <= 0;  @(posedge clock);
												data [0] <= 1;		@(posedge clock);
						   data [1] <= 1; data [0] <= 0;		@(posedge clock);
												data [0] <= 1;		@(posedge clock);
							data [3] <= 1; data [2:0] <= 0;  @(posedge clock);
												data [0] <= 1;		@(posedge clock);
						   data [1] <= 1; data [0] <= 0;		@(posedge clock);
												data [0] <= 1;		@(posedge clock);
							data [2] <= 1;	data [1:0] <= 0;  @(posedge clock);
												data [0] <= 1;		@(posedge clock);
						   data [1] <= 1; data [0] <= 0;		@(posedge clock);
												data [0] <= 1;		@(posedge clock);					
					address [0] <= 1;								@(posedge clock);
							data [0] <= 1;							@(posedge clock);
						   data [1] <= 1; data [0] <= 0;		@(posedge clock);
												data [0] <= 1;		@(posedge clock);
							data [2] <= 1;	data [1:0] <= 0;  @(posedge clock);
												data [0] <= 1;		@(posedge clock);
						   data [1] <= 1; data [0] <= 0;		@(posedge clock);
												data [0] <= 1;		@(posedge clock);
							data [3] <= 1; data [2:0] <= 0;  @(posedge clock);
												data [0] <= 1;		@(posedge clock);
						   data [1] <= 1; data [0] <= 0;		@(posedge clock);
												data [0] <= 1;		@(posedge clock);
							data [2] <= 1;	data [1:0] <= 0;  @(posedge clock);
												data [0] <= 1;		@(posedge clock);
						   data [1] <= 1; data [0] <= 0;		@(posedge clock);
												data [0] <= 1;		@(posedge clock);					
					address [3] <= 1; address [2:0] <= 0;  @(posedge clock);
							data [0] <= 1;							@(posedge clock);
						   data [1] <= 1; data [0] <= 0;		@(posedge clock);
												data [0] <= 1;		@(posedge clock);
							data [2] <= 1;	data [1:0] <= 0;  @(posedge clock);
												data [0] <= 1;		@(posedge clock);
						   data [1] <= 1; data [0] <= 0;		@(posedge clock);
												data [0] <= 1;		@(posedge clock);
							data [3] <= 1; data [2:0] <= 0;  @(posedge clock);
												data [0] <= 1;		@(posedge clock);
						   data [1] <= 1; data [0] <= 0;		@(posedge clock);
												data [0] <= 1;		@(posedge clock);
							data [2] <= 1;	data [1:0] <= 0;  @(posedge clock);
												data [0] <= 1;		@(posedge clock);
						   data [1] <= 1; data [0] <= 0;		@(posedge clock);
												data [0] <= 1;		@(posedge clock);					
					address [0] <= 1;								@(posedge clock);
							data [0] <= 1;							@(posedge clock);
						   data [1] <= 1; data [0] <= 0;		@(posedge clock);
												data [0] <= 1;		@(posedge clock);
							data [2] <= 1;	data [1:0] <= 0;  @(posedge clock);
												data [0] <= 1;		@(posedge clock);
						   data [1] <= 1; data [0] <= 0;		@(posedge clock);
												data [0] <= 1;		@(posedge clock);
							data [3] <= 1; data [2:0] <= 0;  @(posedge clock);
												data [0] <= 1;		@(posedge clock);
						   data [1] <= 1; data [0] <= 0;		@(posedge clock);
												data [0] <= 1;		@(posedge clock);
							data [2] <= 1;	data [1:0] <= 0;  @(posedge clock);
												data [0] <= 1;		@(posedge clock);
						   data [1] <= 1; data [0] <= 0;		@(posedge clock);
												data [0] <= 1;		@(posedge clock);					
					address [1] <= 1; address [0] <= 0;		@(posedge clock);
							data [0] <= 1;							@(posedge clock);
						   data [1] <= 1; data [0] <= 0;		@(posedge clock);
												data [0] <= 1;		@(posedge clock);
							data [2] <= 1;	data [1:0] <= 0;  @(posedge clock);
												data [0] <= 1;		@(posedge clock);
						   data [1] <= 1; data [0] <= 0;		@(posedge clock);
												data [0] <= 1;		@(posedge clock);
							data [3] <= 1; data [2:0] <= 0;  @(posedge clock);
												data [0] <= 1;		@(posedge clock);
						   data [1] <= 1; data [0] <= 0;		@(posedge clock);
												data [0] <= 1;		@(posedge clock);
							data [2] <= 1;	data [1:0] <= 0;  @(posedge clock);
												data [0] <= 1;		@(posedge clock);
						   data [1] <= 1; data [0] <= 0;		@(posedge clock);
												data [0] <= 1;		@(posedge clock);					
					address [0] <= 1;								@(posedge clock);
							data [0] <= 1;							@(posedge clock);
						   data [1] <= 1; data [0] <= 0;		@(posedge clock);
												data [0] <= 1;		@(posedge clock);
							data [2] <= 1;	data [1:0] <= 0;  @(posedge clock);
												data [0] <= 1;		@(posedge clock);
						   data [1] <= 1; data [0] <= 0;		@(posedge clock);
												data [0] <= 1;		@(posedge clock);
							data [3] <= 1; data [2:0] <= 0;  @(posedge clock);
												data [0] <= 1;		@(posedge clock);
						   data [1] <= 1; data [0] <= 0;		@(posedge clock);
												data [0] <= 1;		@(posedge clock);
							data [2] <= 1;	data [1:0] <= 0;  @(posedge clock);
												data [0] <= 1;		@(posedge clock);
						   data [1] <= 1; data [0] <= 0;		@(posedge clock);
												data [0] <= 1;		@(posedge clock);					
					address [2] <= 1; address [1:0] <= 0;  @(posedge clock);
							data [0] <= 1;							@(posedge clock);
						   data [1] <= 1; data [0] <= 0;		@(posedge clock);
												data [0] <= 1;		@(posedge clock);
							data [2] <= 1;	data [1:0] <= 0;  @(posedge clock);
												data [0] <= 1;		@(posedge clock);
						   data [1] <= 1; data [0] <= 0;		@(posedge clock);
												data [0] <= 1;		@(posedge clock);
							data [3] <= 1; data [2:0] <= 0;  @(posedge clock);
												data [0] <= 1;		@(posedge clock);
						   data [1] <= 1; data [0] <= 0;		@(posedge clock);
												data [0] <= 1;		@(posedge clock);
							data [2] <= 1;	data [1:0] <= 0;  @(posedge clock);
												data [0] <= 1;		@(posedge clock);
						   data [1] <= 1; data [0] <= 0;		@(posedge clock);
												data [0] <= 1;		@(posedge clock);					
					address [0] <= 1; 							@(posedge clock);
							data [0] <= 1;							@(posedge clock);
						   data [1] <= 1; data [0] <= 0;		@(posedge clock);
												data [0] <= 1;		@(posedge clock);
							data [2] <= 1;	data [1:0] <= 0;  @(posedge clock);
												data [0] <= 1;		@(posedge clock);
						   data [1] <= 1; data [0] <= 0;		@(posedge clock);
												data [0] <= 1;		@(posedge clock);
							data [3] <= 1; data [2:0] <= 0;  @(posedge clock);
												data [0] <= 1;		@(posedge clock);
						   data [1] <= 1; data [0] <= 0;		@(posedge clock);
												data [0] <= 1;		@(posedge clock);
							data [2] <= 1;	data [1:0] <= 0;  @(posedge clock);
												data [0] <= 1;		@(posedge clock);
						   data [1] <= 1; data [0] <= 0;		@(posedge clock);
												data [0] <= 1;		@(posedge clock);					
					address [1] <= 1; address [0] <= 0;    @(posedge clock);
							data [0] <= 1;							@(posedge clock);
						   data [1] <= 1; data [0] <= 0;		@(posedge clock);
												data [0] <= 1;		@(posedge clock);
							data [2] <= 1;	data [1:0] <= 0;  @(posedge clock);
												data [0] <= 1;		@(posedge clock);
						   data [1] <= 1; data [0] <= 0;		@(posedge clock);
												data [0] <= 1;		@(posedge clock);
							data [3] <= 1; data [2:0] <= 0;  @(posedge clock);
												data [0] <= 1;		@(posedge clock);
						   data [1] <= 1; data [0] <= 0;		@(posedge clock);
												data [0] <= 1;		@(posedge clock);
							data [2] <= 1;	data [1:0] <= 0;  @(posedge clock);
												data [0] <= 1;		@(posedge clock);
						   data [1] <= 1; data [0] <= 0;		@(posedge clock);
												data [0] <= 1;		@(posedge clock);					
					address [0] <= 1;								@(posedge clock);
							data [0] <= 1;							@(posedge clock);
						   data [1] <= 1; data [0] <= 0;		@(posedge clock);
												data [0] <= 1;		@(posedge clock);
							data [2] <= 1;	data [1:0] <= 0;  @(posedge clock);
												data [0] <= 1;		@(posedge clock);
						   data [1] <= 1; data [0] <= 0;		@(posedge clock);
												data [0] <= 1;		@(posedge clock);
							data [3] <= 1; data [2:0] <= 0;  @(posedge clock);
												data [0] <= 1;		@(posedge clock);
						   data [1] <= 1; data [0] <= 0;		@(posedge clock);
												data [0] <= 1;		@(posedge clock);
							data [2] <= 1;	data [1:0] <= 0;  @(posedge clock);
												data [0] <= 1;		@(posedge clock);
						   data [1] <= 1; data [0] <= 0;		@(posedge clock);
												data [0] <= 1;		@(posedge clock);					
					address [4] <= 1;	address [3:0] <= 0;	@(posedge clock);
							data [0] <= 1;							@(posedge clock);
						   data [1] <= 1; data [0] <= 0;		@(posedge clock);
												data [0] <= 1;		@(posedge clock);
							data [2] <= 1;	data [1:0] <= 0;  @(posedge clock);
												data [0] <= 1;		@(posedge clock);
						   data [1] <= 1; data [0] <= 0;		@(posedge clock);
												data [0] <= 1;		@(posedge clock);
							data [3] <= 1; data [2:0] <= 0;  @(posedge clock);
												data [0] <= 1;		@(posedge clock);
						   data [1] <= 1; data [0] <= 0;		@(posedge clock);
												data [0] <= 1;		@(posedge clock);
							data [2] <= 1;	data [1:0] <= 0;  @(posedge clock);
												data [0] <= 1;		@(posedge clock);
						   data [1] <= 1; data [0] <= 0;		@(posedge clock);
												data [0] <= 1;		@(posedge clock);					
					address [0] <= 1;								@(posedge clock); 
							data [0] <= 1;							@(posedge clock);
						   data [1] <= 1; data [0] <= 0;		@(posedge clock);
												data [0] <= 1;		@(posedge clock);
							data [2] <= 1;	data [1:0] <= 0;  @(posedge clock);
												data [0] <= 1;		@(posedge clock);
						   data [1] <= 1; data [0] <= 0;		@(posedge clock);
												data [0] <= 1;		@(posedge clock);
							data [3] <= 1; data [2:0] <= 0;  @(posedge clock);
												data [0] <= 1;		@(posedge clock);
						   data [1] <= 1; data [0] <= 0;		@(posedge clock);
												data [0] <= 1;		@(posedge clock);
							data [2] <= 1;	data [1:0] <= 0;  @(posedge clock);
												data [0] <= 1;		@(posedge clock);
						   data [1] <= 1; data [0] <= 0;		@(posedge clock);
												data [0] <= 1;		@(posedge clock);					
					address [1] <= 1; address [0] <= 0;		@(posedge clock);
							data [0] <= 1;							@(posedge clock);
						   data [1] <= 1; data [0] <= 0;		@(posedge clock);
												data [0] <= 1;		@(posedge clock);
							data [2] <= 1;	data [1:0] <= 0;  @(posedge clock);
												data [0] <= 1;		@(posedge clock);
						   data [1] <= 1; data [0] <= 0;		@(posedge clock);
												data [0] <= 1;		@(posedge clock);
							data [3] <= 1; data [2:0] <= 0;  @(posedge clock);
												data [0] <= 1;		@(posedge clock);
						   data [1] <= 1; data [0] <= 0;		@(posedge clock);
												data [0] <= 1;		@(posedge clock);
							data [2] <= 1;	data [1:0] <= 0;  @(posedge clock);
												data [0] <= 1;		@(posedge clock);
						   data [1] <= 1; data [0] <= 0;		@(posedge clock);
												data [0] <= 1;		@(posedge clock);					
					address [0] <= 1;								@(posedge clock);
							data [0] <= 1;							@(posedge clock);
						   data [1] <= 1; data [0] <= 0;		@(posedge clock);
												data [0] <= 1;		@(posedge clock);
							data [2] <= 1;	data [1:0] <= 0;  @(posedge clock);
												data [0] <= 1;		@(posedge clock);
						   data [1] <= 1; data [0] <= 0;		@(posedge clock);
												data [0] <= 1;		@(posedge clock);
							data [3] <= 1; data [2:0] <= 0;  @(posedge clock);
												data [0] <= 1;		@(posedge clock);
						   data [1] <= 1; data [0] <= 0;		@(posedge clock);
												data [0] <= 1;		@(posedge clock);
							data [2] <= 1;	data [1:0] <= 0;  @(posedge clock);
												data [0] <= 1;		@(posedge clock);
						   data [1] <= 1; data [0] <= 0;		@(posedge clock);
												data [0] <= 1;		@(posedge clock);					
					address [2] <= 1; address [1:0] <= 0;  @(posedge clock);
							data [0] <= 1;							@(posedge clock);
						   data [1] <= 1; data [0] <= 0;		@(posedge clock);
												data [0] <= 1;		@(posedge clock);
							data [2] <= 1;	data [1:0] <= 0;  @(posedge clock);
												data [0] <= 1;		@(posedge clock);
						   data [1] <= 1; data [0] <= 0;		@(posedge clock);
												data [0] <= 1;		@(posedge clock);
							data [3] <= 1; data [2:0] <= 0;  @(posedge clock);
												data [0] <= 1;		@(posedge clock);
						   data [1] <= 1; data [0] <= 0;		@(posedge clock);
												data [0] <= 1;		@(posedge clock);
							data [2] <= 1;	data [1:0] <= 0;  @(posedge clock);
												data [0] <= 1;		@(posedge clock);
						   data [1] <= 1; data [0] <= 0;		@(posedge clock);
												data [0] <= 1;		@(posedge clock);					
					address [0] <= 1; 							@(posedge clock);
							data [0] <= 1;							@(posedge clock);
						   data [1] <= 1; data [0] <= 0;		@(posedge clock);
												data [0] <= 1;		@(posedge clock);
							data [2] <= 1;	data [1:0] <= 0;  @(posedge clock);
												data [0] <= 1;		@(posedge clock);
						   data [1] <= 1; data [0] <= 0;		@(posedge clock);
												data [0] <= 1;		@(posedge clock);
							data [3] <= 1; data [2:0] <= 0;  @(posedge clock);
												data [0] <= 1;		@(posedge clock);
						   data [1] <= 1; data [0] <= 0;		@(posedge clock);
												data [0] <= 1;		@(posedge clock);
							data [2] <= 1;	data [1:0] <= 0;  @(posedge clock);
												data [0] <= 1;		@(posedge clock);
						   data [1] <= 1; data [0] <= 0;		@(posedge clock);
												data [0] <= 1;		@(posedge clock);					
					address [1] <= 1; address [0] <= 0;    @(posedge clock);
							data [0] <= 1;							@(posedge clock);
						   data [1] <= 1; data [0] <= 0;		@(posedge clock);
												data [0] <= 1;		@(posedge clock);
							data [2] <= 1;	data [1:0] <= 0;  @(posedge clock);
												data [0] <= 1;		@(posedge clock);
						   data [1] <= 1; data [0] <= 0;		@(posedge clock);
												data [0] <= 1;		@(posedge clock);
							data [3] <= 1; data [2:0] <= 0;  @(posedge clock);
												data [0] <= 1;		@(posedge clock);
						   data [1] <= 1; data [0] <= 0;		@(posedge clock);
												data [0] <= 1;		@(posedge clock);
							data [2] <= 1;	data [1:0] <= 0;  @(posedge clock);
												data [0] <= 1;		@(posedge clock);
						   data [1] <= 1; data [0] <= 0;		@(posedge clock);
												data [0] <= 1;		@(posedge clock);					
					address [0] <= 1;								@(posedge clock);
							data [0] <= 1;							@(posedge clock);
						   data [1] <= 1; data [0] <= 0;		@(posedge clock);
												data [0] <= 1;		@(posedge clock);
							data [2] <= 1;	data [1:0] <= 0;  @(posedge clock);
												data [0] <= 1;		@(posedge clock);
						   data [1] <= 1; data [0] <= 0;		@(posedge clock);
												data [0] <= 1;		@(posedge clock);
							data [3] <= 1; data [2:0] <= 0;  @(posedge clock);
												data [0] <= 1;		@(posedge clock);
						   data [1] <= 1; data [0] <= 0;		@(posedge clock);
												data [0] <= 1;		@(posedge clock);
							data [2] <= 1;	data [1:0] <= 0;  @(posedge clock);
												data [0] <= 1;		@(posedge clock);
						   data [1] <= 1; data [0] <= 0;		@(posedge clock);
												data [0] <= 1;		@(posedge clock);					
					address [3] <= 1; address [2:0] <= 0;  @(posedge clock);
							data [0] <= 1;							@(posedge clock);
						   data [1] <= 1; data [0] <= 0;		@(posedge clock);
												data [0] <= 1;		@(posedge clock);
							data [2] <= 1;	data [1:0] <= 0;  @(posedge clock);
												data [0] <= 1;		@(posedge clock);
						   data [1] <= 1; data [0] <= 0;		@(posedge clock);
												data [0] <= 1;		@(posedge clock);
							data [3] <= 1; data [2:0] <= 0;  @(posedge clock);
												data [0] <= 1;		@(posedge clock);
						   data [1] <= 1; data [0] <= 0;		@(posedge clock);
												data [0] <= 1;		@(posedge clock);
							data [2] <= 1;	data [1:0] <= 0;  @(posedge clock);
												data [0] <= 1;		@(posedge clock);
						   data [1] <= 1; data [0] <= 0;		@(posedge clock);
												data [0] <= 1;		@(posedge clock);					
					address [0] <= 1;								@(posedge clock);
							data [0] <= 1;							@(posedge clock);
						   data [1] <= 1; data [0] <= 0;		@(posedge clock);
												data [0] <= 1;		@(posedge clock);
							data [2] <= 1;	data [1:0] <= 0;  @(posedge clock);
												data [0] <= 1;		@(posedge clock);
						   data [1] <= 1; data [0] <= 0;		@(posedge clock);
												data [0] <= 1;		@(posedge clock);
							data [3] <= 1; data [2:0] <= 0;  @(posedge clock);
												data [0] <= 1;		@(posedge clock);
						   data [1] <= 1; data [0] <= 0;		@(posedge clock);
												data [0] <= 1;		@(posedge clock);
							data [2] <= 1;	data [1:0] <= 0;  @(posedge clock);
												data [0] <= 1;		@(posedge clock);
						   data [1] <= 1; data [0] <= 0;		@(posedge clock);
												data [0] <= 1;		@(posedge clock);					
					address [1] <= 1; address [0] <= 0;		@(posedge clock);
							data [0] <= 1;							@(posedge clock);
						   data [1] <= 1; data [0] <= 0;		@(posedge clock);
												data [0] <= 1;		@(posedge clock);
							data [2] <= 1;	data [1:0] <= 0;  @(posedge clock);
												data [0] <= 1;		@(posedge clock);
						   data [1] <= 1; data [0] <= 0;		@(posedge clock);
												data [0] <= 1;		@(posedge clock);
							data [3] <= 1; data [2:0] <= 0;  @(posedge clock);
												data [0] <= 1;		@(posedge clock);
						   data [1] <= 1; data [0] <= 0;		@(posedge clock);
												data [0] <= 1;		@(posedge clock);
							data [2] <= 1;	data [1:0] <= 0;  @(posedge clock);
												data [0] <= 1;		@(posedge clock);
						   data [1] <= 1; data [0] <= 0;		@(posedge clock);
												data [0] <= 1;		@(posedge clock);					
					address [0] <= 1;								@(posedge clock);
							data [0] <= 1;							@(posedge clock);
						   data [1] <= 1; data [0] <= 0;		@(posedge clock);
												data [0] <= 1;		@(posedge clock);
							data [2] <= 1;	data [1:0] <= 0;  @(posedge clock);
												data [0] <= 1;		@(posedge clock);
						   data [1] <= 1; data [0] <= 0;		@(posedge clock);
												data [0] <= 1;		@(posedge clock);
							data [3] <= 1; data [2:0] <= 0;  @(posedge clock);
												data [0] <= 1;		@(posedge clock);
						   data [1] <= 1; data [0] <= 0;		@(posedge clock);
												data [0] <= 1;		@(posedge clock);
							data [2] <= 1;	data [1:0] <= 0;  @(posedge clock);
												data [0] <= 1;		@(posedge clock);
						   data [1] <= 1; data [0] <= 0;		@(posedge clock);
												data [0] <= 1;		@(posedge clock);					
					address [2] <= 1; address [1:0] <= 0;  @(posedge clock);
							data [0] <= 1;							@(posedge clock);
						   data [1] <= 1; data [0] <= 0;		@(posedge clock);
												data [0] <= 1;		@(posedge clock);
							data [2] <= 1;	data [1:0] <= 0;  @(posedge clock);
												data [0] <= 1;		@(posedge clock);
						   data [1] <= 1; data [0] <= 0;		@(posedge clock);
												data [0] <= 1;		@(posedge clock);
							data [3] <= 1; data [2:0] <= 0;  @(posedge clock);
												data [0] <= 1;		@(posedge clock);
						   data [1] <= 1; data [0] <= 0;		@(posedge clock);
												data [0] <= 1;		@(posedge clock);
							data [2] <= 1;	data [1:0] <= 0;  @(posedge clock);
												data [0] <= 1;		@(posedge clock);
						   data [1] <= 1; data [0] <= 0;		@(posedge clock);
												data [0] <= 1;		@(posedge clock);					
					address [0] <= 1; 							@(posedge clock);
							data [0] <= 1;							@(posedge clock);
						   data [1] <= 1; data [0] <= 0;		@(posedge clock);
												data [0] <= 1;		@(posedge clock);
							data [2] <= 1;	data [1:0] <= 0;  @(posedge clock);
												data [0] <= 1;		@(posedge clock);
						   data [1] <= 1; data [0] <= 0;		@(posedge clock);
												data [0] <= 1;		@(posedge clock);
							data [3] <= 1; data [2:0] <= 0;  @(posedge clock);
												data [0] <= 1;		@(posedge clock);
						   data [1] <= 1; data [0] <= 0;		@(posedge clock);
												data [0] <= 1;		@(posedge clock);
							data [2] <= 1;	data [1:0] <= 0;  @(posedge clock);
												data [0] <= 1;		@(posedge clock);
						   data [1] <= 1; data [0] <= 0;		@(posedge clock);
												data [0] <= 1;		@(posedge clock);					
					address [1] <= 1; address [0] <= 0;    @(posedge clock);
							data [0] <= 1;							@(posedge clock);
						   data [1] <= 1; data [0] <= 0;		@(posedge clock);
												data [0] <= 1;		@(posedge clock);
							data [2] <= 1;	data [1:0] <= 0;  @(posedge clock);
												data [0] <= 1;		@(posedge clock);
						   data [1] <= 1; data [0] <= 0;		@(posedge clock);
												data [0] <= 1;		@(posedge clock);
							data [3] <= 1; data [2:0] <= 0;  @(posedge clock);
												data [0] <= 1;		@(posedge clock);
						   data [1] <= 1; data [0] <= 0;		@(posedge clock);
												data [0] <= 1;		@(posedge clock);
							data [2] <= 1;	data [1:0] <= 0;  @(posedge clock);
												data [0] <= 1;		@(posedge clock);
						   data [1] <= 1; data [0] <= 0;		@(posedge clock);
												data [0] <= 1;		@(posedge clock);					
					address [0] <= 1;								@(posedge clock);
							data [0] <= 1;							@(posedge clock);
						   data [1] <= 1; data [0] <= 0;		@(posedge clock);
												data [0] <= 1;		@(posedge clock);
							data [2] <= 1;	data [1:0] <= 0;  @(posedge clock);
												data [0] <= 1;		@(posedge clock);
						   data [1] <= 1; data [0] <= 0;		@(posedge clock);
												data [0] <= 1;		@(posedge clock);
							data [3] <= 1; data [2:0] <= 0;  @(posedge clock);
												data [0] <= 1;		@(posedge clock);
						   data [1] <= 1; data [0] <= 0;		@(posedge clock);
												data [0] <= 1;		@(posedge clock);
							data [2] <= 1;	data [1:0] <= 0;  @(posedge clock);
												data [0] <= 1;		@(posedge clock);
						   data [1] <= 1; data [0] <= 0;		@(posedge clock);
												data [0] <= 1;		@(posedge clock);
																								// do it all again
	wren <= 1;  address [4:0] <= 0;  data [2:0] <= 0;  @(posedge clock);
												data [0] <= 1;		@(posedge clock);
						   data [1] <= 1; data [0] <= 0;		@(posedge clock);
												data [0] <= 1;		@(posedge clock);
							data [2] <= 1;	data [1:0] <= 0;  @(posedge clock);
												data [0] <= 1;		@(posedge clock);
						   data [1] <= 1; data [0] <= 0;		@(posedge clock);
												data [0] <= 1;		@(posedge clock);
							data [3] <= 1; data [2:0] <= 0;  @(posedge clock);
												data [0] <= 1;		@(posedge clock);
						   data [1] <= 1; data [0] <= 0;		@(posedge clock);
												data [0] <= 1;		@(posedge clock);
							data [2] <= 1;	data [1:0] <= 0;  @(posedge clock);
												data [0] <= 1;		@(posedge clock);
						   data [1] <= 1; data [0] <= 0;		@(posedge clock);
												data [0] <= 1;		@(posedge clock);
					address [0] <= 1;								@(posedge clock);
							data [0] <= 1;							@(posedge clock);
						   data [1] <= 1; data [0] <= 0;		@(posedge clock);
												data [0] <= 1;		@(posedge clock);
							data [2] <= 1;	data [1:0] <= 0;  @(posedge clock);
												data [0] <= 1;		@(posedge clock);
						   data [1] <= 1; data [0] <= 0;		@(posedge clock);
												data [0] <= 1;		@(posedge clock);
							data [3] <= 1; data [2:0] <= 0;  @(posedge clock);
												data [0] <= 1;		@(posedge clock);
						   data [1] <= 1; data [0] <= 0;		@(posedge clock);
												data [0] <= 1;		@(posedge clock);
							data [2] <= 1;	data [1:0] <= 0;  @(posedge clock);
												data [0] <= 1;		@(posedge clock);
						   data [1] <= 1; data [0] <= 0;		@(posedge clock);
												data [0] <= 1;		@(posedge clock);
					address [1] <= 1; address [0] <= 0;		@(posedge clock);
							data [0] <= 1;							@(posedge clock);
						   data [1] <= 1; data [0] <= 0;		@(posedge clock);
												data [0] <= 1;		@(posedge clock);
							data [2] <= 1;	data [1:0] <= 0;  @(posedge clock);
												data [0] <= 1;		@(posedge clock);
						   data [1] <= 1; data [0] <= 0;		@(posedge clock);
												data [0] <= 1;		@(posedge clock);
							data [3] <= 1; data [2:0] <= 0;  @(posedge clock);
												data [0] <= 1;		@(posedge clock);
						   data [1] <= 1; data [0] <= 0;		@(posedge clock);
												data [0] <= 1;		@(posedge clock);
							data [2] <= 1;	data [1:0] <= 0;  @(posedge clock);
												data [0] <= 1;		@(posedge clock);
						   data [1] <= 1; data [0] <= 0;		@(posedge clock);
												data [0] <= 1;		@(posedge clock);					
					address [0] <= 1;								@(posedge clock);
							data [0] <= 1;							@(posedge clock);
						   data [1] <= 1; data [0] <= 0;		@(posedge clock);
												data [0] <= 1;		@(posedge clock);
							data [2] <= 1;	data [1:0] <= 0;  @(posedge clock);
												data [0] <= 1;		@(posedge clock);
						   data [1] <= 1; data [0] <= 0;		@(posedge clock);
												data [0] <= 1;		@(posedge clock);
							data [3] <= 1; data [2:0] <= 0;  @(posedge clock);
												data [0] <= 1;		@(posedge clock);
						   data [1] <= 1; data [0] <= 0;		@(posedge clock);
												data [0] <= 1;		@(posedge clock);
							data [2] <= 1;	data [1:0] <= 0;  @(posedge clock);
												data [0] <= 1;		@(posedge clock);
						   data [1] <= 1; data [0] <= 0;		@(posedge clock);
												data [0] <= 1;		@(posedge clock);					
					address [2] <= 1; address [1:0] <= 0;  @(posedge clock);
							data [0] <= 1;							@(posedge clock);
						   data [1] <= 1; data [0] <= 0;		@(posedge clock);
												data [0] <= 1;		@(posedge clock);
							data [2] <= 1;	data [1:0] <= 0;  @(posedge clock);
												data [0] <= 1;		@(posedge clock);
						   data [1] <= 1; data [0] <= 0;		@(posedge clock);
												data [0] <= 1;		@(posedge clock);
							data [3] <= 1; data [2:0] <= 0;  @(posedge clock);
												data [0] <= 1;		@(posedge clock);
						   data [1] <= 1; data [0] <= 0;		@(posedge clock);
												data [0] <= 1;		@(posedge clock);
							data [2] <= 1;	data [1:0] <= 0;  @(posedge clock);
												data [0] <= 1;		@(posedge clock);
						   data [1] <= 1; data [0] <= 0;		@(posedge clock);
												data [0] <= 1;		@(posedge clock);					
					address [0] <= 1; 							@(posedge clock);
							data [0] <= 1;							@(posedge clock);
						   data [1] <= 1; data [0] <= 0;		@(posedge clock);
												data [0] <= 1;		@(posedge clock);
							data [2] <= 1;	data [1:0] <= 0;  @(posedge clock);
												data [0] <= 1;		@(posedge clock);
						   data [1] <= 1; data [0] <= 0;		@(posedge clock);
												data [0] <= 1;		@(posedge clock);
							data [3] <= 1; data [2:0] <= 0;  @(posedge clock);
												data [0] <= 1;		@(posedge clock);
						   data [1] <= 1; data [0] <= 0;		@(posedge clock);
												data [0] <= 1;		@(posedge clock);
							data [2] <= 1;	data [1:0] <= 0;  @(posedge clock);
												data [0] <= 1;		@(posedge clock);
						   data [1] <= 1; data [0] <= 0;		@(posedge clock);
												data [0] <= 1;		@(posedge clock);					
					address [1] <= 1; address [0] <= 0;    @(posedge clock);
							data [0] <= 1;							@(posedge clock);
						   data [1] <= 1; data [0] <= 0;		@(posedge clock);
												data [0] <= 1;		@(posedge clock);
							data [2] <= 1;	data [1:0] <= 0;  @(posedge clock);
												data [0] <= 1;		@(posedge clock);
						   data [1] <= 1; data [0] <= 0;		@(posedge clock);
												data [0] <= 1;		@(posedge clock);
							data [3] <= 1; data [2:0] <= 0;  @(posedge clock);
												data [0] <= 1;		@(posedge clock);
						   data [1] <= 1; data [0] <= 0;		@(posedge clock);
												data [0] <= 1;		@(posedge clock);
							data [2] <= 1;	data [1:0] <= 0;  @(posedge clock);
												data [0] <= 1;		@(posedge clock);
						   data [1] <= 1; data [0] <= 0;		@(posedge clock);
												data [0] <= 1;		@(posedge clock);					
					address [0] <= 1;								@(posedge clock);
							data [0] <= 1;							@(posedge clock);
						   data [1] <= 1; data [0] <= 0;		@(posedge clock);
												data [0] <= 1;		@(posedge clock);
							data [2] <= 1;	data [1:0] <= 0;  @(posedge clock);
												data [0] <= 1;		@(posedge clock);
						   data [1] <= 1; data [0] <= 0;		@(posedge clock);
												data [0] <= 1;		@(posedge clock);
							data [3] <= 1; data [2:0] <= 0;  @(posedge clock);
												data [0] <= 1;		@(posedge clock);
						   data [1] <= 1; data [0] <= 0;		@(posedge clock);
												data [0] <= 1;		@(posedge clock);
							data [2] <= 1;	data [1:0] <= 0;  @(posedge clock);
												data [0] <= 1;		@(posedge clock);
						   data [1] <= 1; data [0] <= 0;		@(posedge clock);
												data [0] <= 1;		@(posedge clock);					
					address [3] <= 1; address [2:0] <= 0;  @(posedge clock);
							data [0] <= 1;							@(posedge clock);
						   data [1] <= 1; data [0] <= 0;		@(posedge clock);
												data [0] <= 1;		@(posedge clock);
							data [2] <= 1;	data [1:0] <= 0;  @(posedge clock);
												data [0] <= 1;		@(posedge clock);
						   data [1] <= 1; data [0] <= 0;		@(posedge clock);
												data [0] <= 1;		@(posedge clock);
							data [3] <= 1; data [2:0] <= 0;  @(posedge clock);
												data [0] <= 1;		@(posedge clock);
						   data [1] <= 1; data [0] <= 0;		@(posedge clock);
												data [0] <= 1;		@(posedge clock);
							data [2] <= 1;	data [1:0] <= 0;  @(posedge clock);
												data [0] <= 1;		@(posedge clock);
						   data [1] <= 1; data [0] <= 0;		@(posedge clock);
												data [0] <= 1;		@(posedge clock);					
					address [0] <= 1;								@(posedge clock);
							data [0] <= 1;							@(posedge clock);
						   data [1] <= 1; data [0] <= 0;		@(posedge clock);
												data [0] <= 1;		@(posedge clock);
							data [2] <= 1;	data [1:0] <= 0;  @(posedge clock);
												data [0] <= 1;		@(posedge clock);
						   data [1] <= 1; data [0] <= 0;		@(posedge clock);
												data [0] <= 1;		@(posedge clock);
							data [3] <= 1; data [2:0] <= 0;  @(posedge clock);
												data [0] <= 1;		@(posedge clock);
						   data [1] <= 1; data [0] <= 0;		@(posedge clock);
												data [0] <= 1;		@(posedge clock);
							data [2] <= 1;	data [1:0] <= 0;  @(posedge clock);
												data [0] <= 1;		@(posedge clock);
						   data [1] <= 1; data [0] <= 0;		@(posedge clock);
												data [0] <= 1;		@(posedge clock);					
					address [1] <= 1; address [0] <= 0;		@(posedge clock);
							data [0] <= 1;							@(posedge clock);
						   data [1] <= 1; data [0] <= 0;		@(posedge clock);
												data [0] <= 1;		@(posedge clock);
							data [2] <= 1;	data [1:0] <= 0;  @(posedge clock);
												data [0] <= 1;		@(posedge clock);
						   data [1] <= 1; data [0] <= 0;		@(posedge clock);
												data [0] <= 1;		@(posedge clock);
							data [3] <= 1; data [2:0] <= 0;  @(posedge clock);
												data [0] <= 1;		@(posedge clock);
						   data [1] <= 1; data [0] <= 0;		@(posedge clock);
												data [0] <= 1;		@(posedge clock);
							data [2] <= 1;	data [1:0] <= 0;  @(posedge clock);
												data [0] <= 1;		@(posedge clock);
						   data [1] <= 1; data [0] <= 0;		@(posedge clock);
												data [0] <= 1;		@(posedge clock);					
					address [0] <= 1;								@(posedge clock);
							data [0] <= 1;							@(posedge clock);
						   data [1] <= 1; data [0] <= 0;		@(posedge clock);
												data [0] <= 1;		@(posedge clock);
							data [2] <= 1;	data [1:0] <= 0;  @(posedge clock);
												data [0] <= 1;		@(posedge clock);
						   data [1] <= 1; data [0] <= 0;		@(posedge clock);
												data [0] <= 1;		@(posedge clock);
							data [3] <= 1; data [2:0] <= 0;  @(posedge clock);
												data [0] <= 1;		@(posedge clock);
						   data [1] <= 1; data [0] <= 0;		@(posedge clock);
												data [0] <= 1;		@(posedge clock);
							data [2] <= 1;	data [1:0] <= 0;  @(posedge clock);
												data [0] <= 1;		@(posedge clock);
						   data [1] <= 1; data [0] <= 0;		@(posedge clock);
												data [0] <= 1;		@(posedge clock);					
					address [2] <= 1; address [1:0] <= 0;  @(posedge clock);
							data [0] <= 1;							@(posedge clock);
						   data [1] <= 1; data [0] <= 0;		@(posedge clock);
												data [0] <= 1;		@(posedge clock);
							data [2] <= 1;	data [1:0] <= 0;  @(posedge clock);
												data [0] <= 1;		@(posedge clock);
						   data [1] <= 1; data [0] <= 0;		@(posedge clock);
												data [0] <= 1;		@(posedge clock);
							data [3] <= 1; data [2:0] <= 0;  @(posedge clock);
												data [0] <= 1;		@(posedge clock);
						   data [1] <= 1; data [0] <= 0;		@(posedge clock);
												data [0] <= 1;		@(posedge clock);
							data [2] <= 1;	data [1:0] <= 0;  @(posedge clock);
												data [0] <= 1;		@(posedge clock);
						   data [1] <= 1; data [0] <= 0;		@(posedge clock);
												data [0] <= 1;		@(posedge clock);					
					address [0] <= 1; 							@(posedge clock);
							data [0] <= 1;							@(posedge clock);
						   data [1] <= 1; data [0] <= 0;		@(posedge clock);
												data [0] <= 1;		@(posedge clock);
							data [2] <= 1;	data [1:0] <= 0;  @(posedge clock);
												data [0] <= 1;		@(posedge clock);
						   data [1] <= 1; data [0] <= 0;		@(posedge clock);
												data [0] <= 1;		@(posedge clock);
							data [3] <= 1; data [2:0] <= 0;  @(posedge clock);
												data [0] <= 1;		@(posedge clock);
						   data [1] <= 1; data [0] <= 0;		@(posedge clock);
												data [0] <= 1;		@(posedge clock);
							data [2] <= 1;	data [1:0] <= 0;  @(posedge clock);
												data [0] <= 1;		@(posedge clock);
						   data [1] <= 1; data [0] <= 0;		@(posedge clock);
												data [0] <= 1;		@(posedge clock);					
					address [1] <= 1; address [0] <= 0;    @(posedge clock);
							data [0] <= 1;							@(posedge clock);
						   data [1] <= 1; data [0] <= 0;		@(posedge clock);
												data [0] <= 1;		@(posedge clock);
							data [2] <= 1;	data [1:0] <= 0;  @(posedge clock);
												data [0] <= 1;		@(posedge clock);
						   data [1] <= 1; data [0] <= 0;		@(posedge clock);
												data [0] <= 1;		@(posedge clock);
							data [3] <= 1; data [2:0] <= 0;  @(posedge clock);
												data [0] <= 1;		@(posedge clock);
						   data [1] <= 1; data [0] <= 0;		@(posedge clock);
												data [0] <= 1;		@(posedge clock);
							data [2] <= 1;	data [1:0] <= 0;  @(posedge clock);
												data [0] <= 1;		@(posedge clock);
						   data [1] <= 1; data [0] <= 0;		@(posedge clock);
												data [0] <= 1;		@(posedge clock);					
					address [0] <= 1;								@(posedge clock);
							data [0] <= 1;							@(posedge clock);
						   data [1] <= 1; data [0] <= 0;		@(posedge clock);
												data [0] <= 1;		@(posedge clock);
							data [2] <= 1;	data [1:0] <= 0;  @(posedge clock);
												data [0] <= 1;		@(posedge clock);
						   data [1] <= 1; data [0] <= 0;		@(posedge clock);
												data [0] <= 1;		@(posedge clock);
							data [3] <= 1; data [2:0] <= 0;  @(posedge clock);
												data [0] <= 1;		@(posedge clock);
						   data [1] <= 1; data [0] <= 0;		@(posedge clock);
												data [0] <= 1;		@(posedge clock);
							data [2] <= 1;	data [1:0] <= 0;  @(posedge clock);
												data [0] <= 1;		@(posedge clock);
						   data [1] <= 1; data [0] <= 0;		@(posedge clock);
												data [0] <= 1;		@(posedge clock);					
					address [4] <= 1;	address [3:0] <= 0;	@(posedge clock);
							data [0] <= 1;							@(posedge clock);
						   data [1] <= 1; data [0] <= 0;		@(posedge clock);
												data [0] <= 1;		@(posedge clock);
							data [2] <= 1;	data [1:0] <= 0;  @(posedge clock);
												data [0] <= 1;		@(posedge clock);
						   data [1] <= 1; data [0] <= 0;		@(posedge clock);
												data [0] <= 1;		@(posedge clock);
							data [3] <= 1; data [2:0] <= 0;  @(posedge clock);
												data [0] <= 1;		@(posedge clock);
						   data [1] <= 1; data [0] <= 0;		@(posedge clock);
												data [0] <= 1;		@(posedge clock);
							data [2] <= 1;	data [1:0] <= 0;  @(posedge clock);
												data [0] <= 1;		@(posedge clock);
						   data [1] <= 1; data [0] <= 0;		@(posedge clock);
												data [0] <= 1;		@(posedge clock);					
					address [0] <= 1;								@(posedge clock); 
							data [0] <= 1;							@(posedge clock);
						   data [1] <= 1; data [0] <= 0;		@(posedge clock);
												data [0] <= 1;		@(posedge clock);
							data [2] <= 1;	data [1:0] <= 0;  @(posedge clock);
												data [0] <= 1;		@(posedge clock);
						   data [1] <= 1; data [0] <= 0;		@(posedge clock);
												data [0] <= 1;		@(posedge clock);
							data [3] <= 1; data [2:0] <= 0;  @(posedge clock);
												data [0] <= 1;		@(posedge clock);
						   data [1] <= 1; data [0] <= 0;		@(posedge clock);
												data [0] <= 1;		@(posedge clock);
							data [2] <= 1;	data [1:0] <= 0;  @(posedge clock);
												data [0] <= 1;		@(posedge clock);
						   data [1] <= 1; data [0] <= 0;		@(posedge clock);
												data [0] <= 1;		@(posedge clock);					
					address [1] <= 1; address [0] <= 0;		@(posedge clock);
							data [0] <= 1;							@(posedge clock);
						   data [1] <= 1; data [0] <= 0;		@(posedge clock);
												data [0] <= 1;		@(posedge clock);
							data [2] <= 1;	data [1:0] <= 0;  @(posedge clock);
												data [0] <= 1;		@(posedge clock);
						   data [1] <= 1; data [0] <= 0;		@(posedge clock);
												data [0] <= 1;		@(posedge clock);
							data [3] <= 1; data [2:0] <= 0;  @(posedge clock);
												data [0] <= 1;		@(posedge clock);
						   data [1] <= 1; data [0] <= 0;		@(posedge clock);
												data [0] <= 1;		@(posedge clock);
							data [2] <= 1;	data [1:0] <= 0;  @(posedge clock);
												data [0] <= 1;		@(posedge clock);
						   data [1] <= 1; data [0] <= 0;		@(posedge clock);
												data [0] <= 1;		@(posedge clock);					
					address [0] <= 1;								@(posedge clock);
							data [0] <= 1;							@(posedge clock);
						   data [1] <= 1; data [0] <= 0;		@(posedge clock);
												data [0] <= 1;		@(posedge clock);
							data [2] <= 1;	data [1:0] <= 0;  @(posedge clock);
												data [0] <= 1;		@(posedge clock);
						   data [1] <= 1; data [0] <= 0;		@(posedge clock);
												data [0] <= 1;		@(posedge clock);
							data [3] <= 1; data [2:0] <= 0;  @(posedge clock);
												data [0] <= 1;		@(posedge clock);
						   data [1] <= 1; data [0] <= 0;		@(posedge clock);
												data [0] <= 1;		@(posedge clock);
							data [2] <= 1;	data [1:0] <= 0;  @(posedge clock);
												data [0] <= 1;		@(posedge clock);
						   data [1] <= 1; data [0] <= 0;		@(posedge clock);
												data [0] <= 1;		@(posedge clock);					
					address [2] <= 1; address [1:0] <= 0;  @(posedge clock);
							data [0] <= 1;							@(posedge clock);
						   data [1] <= 1; data [0] <= 0;		@(posedge clock);
												data [0] <= 1;		@(posedge clock);
							data [2] <= 1;	data [1:0] <= 0;  @(posedge clock);
												data [0] <= 1;		@(posedge clock);
						   data [1] <= 1; data [0] <= 0;		@(posedge clock);
												data [0] <= 1;		@(posedge clock);
							data [3] <= 1; data [2:0] <= 0;  @(posedge clock);
												data [0] <= 1;		@(posedge clock);
						   data [1] <= 1; data [0] <= 0;		@(posedge clock);
												data [0] <= 1;		@(posedge clock);
							data [2] <= 1;	data [1:0] <= 0;  @(posedge clock);
												data [0] <= 1;		@(posedge clock);
						   data [1] <= 1; data [0] <= 0;		@(posedge clock);
												data [0] <= 1;		@(posedge clock);					
					address [0] <= 1; 							@(posedge clock);
							data [0] <= 1;							@(posedge clock);
						   data [1] <= 1; data [0] <= 0;		@(posedge clock);
												data [0] <= 1;		@(posedge clock);
							data [2] <= 1;	data [1:0] <= 0;  @(posedge clock);
												data [0] <= 1;		@(posedge clock);
						   data [1] <= 1; data [0] <= 0;		@(posedge clock);
												data [0] <= 1;		@(posedge clock);
							data [3] <= 1; data [2:0] <= 0;  @(posedge clock);
												data [0] <= 1;		@(posedge clock);
						   data [1] <= 1; data [0] <= 0;		@(posedge clock);
												data [0] <= 1;		@(posedge clock);
							data [2] <= 1;	data [1:0] <= 0;  @(posedge clock);
												data [0] <= 1;		@(posedge clock);
						   data [1] <= 1; data [0] <= 0;		@(posedge clock);
												data [0] <= 1;		@(posedge clock);					
					address [1] <= 1; address [0] <= 0;    @(posedge clock);
							data [0] <= 1;							@(posedge clock);
						   data [1] <= 1; data [0] <= 0;		@(posedge clock);
												data [0] <= 1;		@(posedge clock);
							data [2] <= 1;	data [1:0] <= 0;  @(posedge clock);
												data [0] <= 1;		@(posedge clock);
						   data [1] <= 1; data [0] <= 0;		@(posedge clock);
												data [0] <= 1;		@(posedge clock);
							data [3] <= 1; data [2:0] <= 0;  @(posedge clock);
												data [0] <= 1;		@(posedge clock);
						   data [1] <= 1; data [0] <= 0;		@(posedge clock);
												data [0] <= 1;		@(posedge clock);
							data [2] <= 1;	data [1:0] <= 0;  @(posedge clock);
												data [0] <= 1;		@(posedge clock);
						   data [1] <= 1; data [0] <= 0;		@(posedge clock);
												data [0] <= 1;		@(posedge clock);					
					address [0] <= 1;								@(posedge clock);
							data [0] <= 1;							@(posedge clock);
						   data [1] <= 1; data [0] <= 0;		@(posedge clock);
												data [0] <= 1;		@(posedge clock);
							data [2] <= 1;	data [1:0] <= 0;  @(posedge clock);
												data [0] <= 1;		@(posedge clock);
						   data [1] <= 1; data [0] <= 0;		@(posedge clock);
												data [0] <= 1;		@(posedge clock);
							data [3] <= 1; data [2:0] <= 0;  @(posedge clock);
												data [0] <= 1;		@(posedge clock);
						   data [1] <= 1; data [0] <= 0;		@(posedge clock);
												data [0] <= 1;		@(posedge clock);
							data [2] <= 1;	data [1:0] <= 0;  @(posedge clock);
												data [0] <= 1;		@(posedge clock);
						   data [1] <= 1; data [0] <= 0;		@(posedge clock);
												data [0] <= 1;		@(posedge clock);					
					address [3] <= 1; address [2:0] <= 0;  @(posedge clock);
							data [0] <= 1;							@(posedge clock);
						   data [1] <= 1; data [0] <= 0;		@(posedge clock);
												data [0] <= 1;		@(posedge clock);
							data [2] <= 1;	data [1:0] <= 0;  @(posedge clock);
												data [0] <= 1;		@(posedge clock);
						   data [1] <= 1; data [0] <= 0;		@(posedge clock);
												data [0] <= 1;		@(posedge clock);
							data [3] <= 1; data [2:0] <= 0;  @(posedge clock);
												data [0] <= 1;		@(posedge clock);
						   data [1] <= 1; data [0] <= 0;		@(posedge clock);
												data [0] <= 1;		@(posedge clock);
							data [2] <= 1;	data [1:0] <= 0;  @(posedge clock);
												data [0] <= 1;		@(posedge clock);
						   data [1] <= 1; data [0] <= 0;		@(posedge clock);
												data [0] <= 1;		@(posedge clock);					
					address [0] <= 1;								@(posedge clock);
							data [0] <= 1;							@(posedge clock);
						   data [1] <= 1; data [0] <= 0;		@(posedge clock);
												data [0] <= 1;		@(posedge clock);
							data [2] <= 1;	data [1:0] <= 0;  @(posedge clock);
												data [0] <= 1;		@(posedge clock);
						   data [1] <= 1; data [0] <= 0;		@(posedge clock);
												data [0] <= 1;		@(posedge clock);
							data [3] <= 1; data [2:0] <= 0;  @(posedge clock);
												data [0] <= 1;		@(posedge clock);
						   data [1] <= 1; data [0] <= 0;		@(posedge clock);
												data [0] <= 1;		@(posedge clock);
							data [2] <= 1;	data [1:0] <= 0;  @(posedge clock);
												data [0] <= 1;		@(posedge clock);
						   data [1] <= 1; data [0] <= 0;		@(posedge clock);
												data [0] <= 1;		@(posedge clock);					
					address [1] <= 1; address [0] <= 0;		@(posedge clock);
							data [0] <= 1;							@(posedge clock);
						   data [1] <= 1; data [0] <= 0;		@(posedge clock);
												data [0] <= 1;		@(posedge clock);
							data [2] <= 1;	data [1:0] <= 0;  @(posedge clock);
												data [0] <= 1;		@(posedge clock);
						   data [1] <= 1; data [0] <= 0;		@(posedge clock);
												data [0] <= 1;		@(posedge clock);
							data [3] <= 1; data [2:0] <= 0;  @(posedge clock);
												data [0] <= 1;		@(posedge clock);
						   data [1] <= 1; data [0] <= 0;		@(posedge clock);
												data [0] <= 1;		@(posedge clock);
							data [2] <= 1;	data [1:0] <= 0;  @(posedge clock);
												data [0] <= 1;		@(posedge clock);
						   data [1] <= 1; data [0] <= 0;		@(posedge clock);
												data [0] <= 1;		@(posedge clock);					
					address [0] <= 1;								@(posedge clock);
							data [0] <= 1;							@(posedge clock);
						   data [1] <= 1; data [0] <= 0;		@(posedge clock);
												data [0] <= 1;		@(posedge clock);
							data [2] <= 1;	data [1:0] <= 0;  @(posedge clock);
												data [0] <= 1;		@(posedge clock);
						   data [1] <= 1; data [0] <= 0;		@(posedge clock);
												data [0] <= 1;		@(posedge clock);
							data [3] <= 1; data [2:0] <= 0;  @(posedge clock);
												data [0] <= 1;		@(posedge clock);
						   data [1] <= 1; data [0] <= 0;		@(posedge clock);
												data [0] <= 1;		@(posedge clock);
							data [2] <= 1;	data [1:0] <= 0;  @(posedge clock);
												data [0] <= 1;		@(posedge clock);
						   data [1] <= 1; data [0] <= 0;		@(posedge clock);
												data [0] <= 1;		@(posedge clock);					
					address [2] <= 1; address [1:0] <= 0;  @(posedge clock);
							data [0] <= 1;							@(posedge clock);
						   data [1] <= 1; data [0] <= 0;		@(posedge clock);
												data [0] <= 1;		@(posedge clock);
							data [2] <= 1;	data [1:0] <= 0;  @(posedge clock);
												data [0] <= 1;		@(posedge clock);
						   data [1] <= 1; data [0] <= 0;		@(posedge clock);
												data [0] <= 1;		@(posedge clock);
							data [3] <= 1; data [2:0] <= 0;  @(posedge clock);
												data [0] <= 1;		@(posedge clock);
						   data [1] <= 1; data [0] <= 0;		@(posedge clock);
												data [0] <= 1;		@(posedge clock);
							data [2] <= 1;	data [1:0] <= 0;  @(posedge clock);
												data [0] <= 1;		@(posedge clock);
						   data [1] <= 1; data [0] <= 0;		@(posedge clock);
												data [0] <= 1;		@(posedge clock);					
					address [0] <= 1; 							@(posedge clock);
							data [0] <= 1;							@(posedge clock);
						   data [1] <= 1; data [0] <= 0;		@(posedge clock);
												data [0] <= 1;		@(posedge clock);
							data [2] <= 1;	data [1:0] <= 0;  @(posedge clock);
												data [0] <= 1;		@(posedge clock);
						   data [1] <= 1; data [0] <= 0;		@(posedge clock);
												data [0] <= 1;		@(posedge clock);
							data [3] <= 1; data [2:0] <= 0;  @(posedge clock);
												data [0] <= 1;		@(posedge clock);
						   data [1] <= 1; data [0] <= 0;		@(posedge clock);
												data [0] <= 1;		@(posedge clock);
							data [2] <= 1;	data [1:0] <= 0;  @(posedge clock);
												data [0] <= 1;		@(posedge clock);
						   data [1] <= 1; data [0] <= 0;		@(posedge clock);
												data [0] <= 1;		@(posedge clock);					
					address [1] <= 1; address [0] <= 0;    @(posedge clock);
							data [0] <= 1;							@(posedge clock);
						   data [1] <= 1; data [0] <= 0;		@(posedge clock);
												data [0] <= 1;		@(posedge clock);
							data [2] <= 1;	data [1:0] <= 0;  @(posedge clock);
												data [0] <= 1;		@(posedge clock);
						   data [1] <= 1; data [0] <= 0;		@(posedge clock);
												data [0] <= 1;		@(posedge clock);
							data [3] <= 1; data [2:0] <= 0;  @(posedge clock);
												data [0] <= 1;		@(posedge clock);
						   data [1] <= 1; data [0] <= 0;		@(posedge clock);
												data [0] <= 1;		@(posedge clock);
							data [2] <= 1;	data [1:0] <= 0;  @(posedge clock);
												data [0] <= 1;		@(posedge clock);
						   data [1] <= 1; data [0] <= 0;		@(posedge clock);
												data [0] <= 1;		@(posedge clock);					
					address [0] <= 1;								@(posedge clock);
							data [0] <= 1;							@(posedge clock);
						   data [1] <= 1; data [0] <= 0;		@(posedge clock);
												data [0] <= 1;		@(posedge clock);
							data [2] <= 1;	data [1:0] <= 0;  @(posedge clock);
												data [0] <= 1;		@(posedge clock);
						   data [1] <= 1; data [0] <= 0;		@(posedge clock);
												data [0] <= 1;		@(posedge clock);
							data [3] <= 1; data [2:0] <= 0;  @(posedge clock);
												data [0] <= 1;		@(posedge clock);
						   data [1] <= 1; data [0] <= 0;		@(posedge clock);
												data [0] <= 1;		@(posedge clock);
							data [2] <= 1;	data [1:0] <= 0;  @(posedge clock);
												data [0] <= 1;		@(posedge clock);
						   data [1] <= 1; data [0] <= 0;		@(posedge clock);
												data [0] <= 1;		@(posedge clock);	
												
	/*wren <= 1;  address [4:0] <= 0;  data [2:0] <= 0;  @(posedge clock);
					address [0] <= 1;								@(posedge clock); 
					address [1] <= 1; address [0] <= 0;		@(posedge clock);
					address [0] <= 1;								@(posedge clock);
					address [2] <= 1; address [1:0] <= 0;  @(posedge clock);
					address [0] <= 1; 							@(posedge clock);
					address [1] <= 1; address [0] <= 0;    @(posedge clock);
					address [0] <= 1;								@(posedge clock);
					address [3] <= 1; address [2:0] <= 0;  @(posedge clock);
					address [0] <= 1;								@(posedge clock);
					address [1] <= 1; address [0] <= 0;		@(posedge clock);
					address [0] <= 1;								@(posedge clock);
					address [2] <= 1; address [1:0] <= 0;  @(posedge clock);
					address [0] <= 1; 							@(posedge clock);
					address [1] <= 1; address [0] <= 0;    @(posedge clock);
					address [0] <= 1;								@(posedge clock);
					address [4] <= 1;	address [3:0] <= 0;	@(posedge clock);
					address [0] <= 1;								@(posedge clock); 
					address [1] <= 1; address [0] <= 0;		@(posedge clock);
					address [0] <= 1;								@(posedge clock);
					address [2] <= 1; address [1:0] <= 0;  @(posedge clock);
					address [0] <= 1; 							@(posedge clock);
					address [1] <= 1; address [0] <= 0;    @(posedge clock);
					address [0] <= 1;								@(posedge clock);
					address [3] <= 1; address [2:0] <= 0;  @(posedge clock);
					address [0] <= 1;								@(posedge clock);
					address [1] <= 1; address [0] <= 0;		@(posedge clock);
					address [0] <= 1;								@(posedge clock);
					address [2] <= 1; address [1:0] <= 0;  @(posedge clock);
					address [0] <= 1; 							@(posedge clock);
					address [1] <= 1; address [0] <= 0;    @(posedge clock);
					address [0] <= 1;								@(posedge clock);
				*/																											
	
	$stop; // End the simulation.  
	end    
endmodule 
	

	